d/inst/Clk5MHz_Clock_clk_wiz_0_0  Jnet (fo=1, routed)X h � ����>��� � � � � � Y
1-Clock_5MHz/ClockingWizzard/inst/clkout1_buf/I  J X h zr�� � � � � � � � r
1-Clock_5MHz/ClockingWizzard/inst/clkout1_buf/OProp_bufg_I_O JBUFGX h zr�����<��� � � � � � M
Segment/CLK  Jnet (fo=11, routed)X h � ��f?��� � � � � � O
#Segment/RefreshCounter_reg[1]/C  JFDREX h zr�� �� � � � � � ��
W  J+(clock Clk5MHz_Clock_clk_wiz_0_0 rise edge)X h zr��    ��� � � � � � :
 Clock_In  J X h zr��    ��� � � � � � `
+'Clock_5MHz/ClockingWizzard/inst/clk_in1  J
net (fo=0)X h � �    ��� � � � � � W
2.Clock_5MHz/ClockingWizzard/inst/clkin1_ibufg/I  J X h � � � � � � � � � s
2.Clock_5MHz/ClockingWizzard/inst/clkin1_ibufg/OProp_ibuf_I_O JIBUFX h zr�����>��� � � � � � z
=9Clock_5MHz/ClockingWizzard/inst/clk_in1_Clock_clk_wiz_0_0  Jnet (fo=1, routed)X h � ����>��� � � � � � ]
84Clock_5MHz/ClockingWizzard/inst/mmcm_adv_inst/CLKIN1  J X h � � � � � � � � � �
95Clock_5MHz/ClockingWizzard/inst/mmcm_adv_inst/CLKOUT0Prop_mmcme2_adv_CLKIN1_CLKOUT0 J
MMCME2_ADVX h zr��C���� � � � � � z
=9Clock_5MHz/ClockingWizzard/inst/Clk5MHz_Cloc